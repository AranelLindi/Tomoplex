----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/25/2023 11:43:05 AM
-- Design Name: 
-- Module Name: SPI_Master_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity SPI_Master_tb is
end;

architecture bench of SPI_Master_tb is
    constant DATA_WIDTH : positive := 8;
    constant Quarz_Taktfrequenz : integer := 100000000;
    constant SPI_Taktfrequenz : integer   :=  20000000;

    component SPI_Master
        Generic ( Quarz_Taktfrequenz : integer;--   := 100000000;
                SPI_Taktfrequenz   : integer;--   :=  30000000;
                DATA_WIDTH             : integer
               );
        Port ( TX_Data  : in  STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
             RX_Data  : out STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
             MOSI     : out STD_LOGIC;
             MISO     : in  STD_LOGIC;
             SCLK     : out STD_LOGIC;
             SS       : out STD_LOGIC;
             TX_Start : in  STD_LOGIC;
             TX_Done  : out STD_LOGIC;
             clk      : in  STD_LOGIC
            );
    end component;

    signal TX_Data: STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0) := (others => '0');
    signal RX_Data: STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
    signal MOSI: STD_LOGIC;
    signal MISO: STD_LOGIC := '0';
    signal SCLK: STD_LOGIC;
    signal SS: STD_LOGIC := '0';
    signal TX_Start: STD_LOGIC := '0';
    signal TX_Done: STD_LOGIC;
    signal clk: STD_LOGIC;

    constant clock_period: time := 10 ns; -- 100 MHz
    -- SPI Clock is generated by DuT and must not necessarily be same value as specified under SPI_Taktfrequenz! So check before implementing it on hardware!
    
    -- Simulates bit stream send process from slave to master.
    -- Because the slave is only allowed to send data when the CS is low a "fake" master transmit process is initiated before and takes place as long as data is written on MISO signal.
    procedure send2Master(constant data : in std_logic_vector(DATA_WIDTH-1 downto 0); signal miso : out std_logic; signal TX_Data : out std_logic_vector(DATA_WIDTH-1 downto 0); signal TX_Start : out std_logic) is
    begin
        wait until rising_edge(CLK);
        
        TX_Data <= (others => '0');
        TX_Start <= '1';
        
        --wait until rising_edge(SCLK);
        for i in data'length-1 downto 0 loop
            wait until rising_edge(SCLK);
            MISO <= data(i);
            
            --wait for SPI_period;
        end loop;       
        
        TX_Start <= '0'; 
    end procedure;
    
    -- Simulates a master transmit process to the slave.
    procedure send2Slave(constant data : in std_logic_vector(DATA_WIDTH-1 downto 0); signal TX_Start : out std_logic; signal TX_Data : out std_logic_vector(DATA_WIDTH-1 downto 0)) is
    begin
        wait until rising_edge(CLK);
        
        TX_Data <= data;
        TX_Start <= '1';
        wait until rising_edge(CLK) and TX_Done = '1';
        TX_Start <= '0';
    end procedure;
begin

    -- Insert values for generic parameters !!
    uut: SPI_Master generic map ( Quarz_Taktfrequenz => Quarz_Taktfrequenz,
                    SPI_Taktfrequenz   => SPI_Taktfrequenz,
                    DATA_WIDTH             => DATA_WIDTH)
        port map ( TX_Data            => TX_Data,
                 RX_Data            => RX_Data,
                 MOSI               => MOSI,
                 MISO               => MISO,
                 SCLK               => SCLK,
                 SS                 => SS,
                 TX_Start           => TX_Start,
                 TX_Done            => TX_Done,
                 clk                => clk );

    stimulus: process
    begin

        -- Put initialisation code here
        wait for 200 ns;
        
        -- Put test bench stimulus code here
        
        -- Send data to master.
        send2Master("10101010", MISO, TX_Data, TX_Start);                
        wait for 200 ns;

        -- Send data from the master to the slave.       
        send2Slave(x"ff", TX_Start, TX_Data);
        wait for 100 ns;
        
        wait;
    end process;

    clocking: process
    begin
        CLK <= '0', '1' after clock_period / 2;
        wait for clock_period;
    end process;
end;